module mynot(
	input in,
	output out
);

	mynand(in, in, out);

endmodule
