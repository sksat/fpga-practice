module top(
	input wire RST_N,
	output wire R_LED
);

assign R_LED = RST_N;

endmodule
